
//`define CONFIG_1 10'b0011111010
//`define CONFIG_2 10'b1100000101
//`define CONFIG_3 10'b1010101010
//`define CONFIG_4 10'b1010101010
//`define CONFIG_5 10'b1011010101
//`define CONFIG_6 10'b0100100101

//`define DATA_1 10'b1010110001
//`define DATA_2 10'b0101001110

//`define ERROR_PROPAGATE_1 10'b0111101000 
//`define ERROR_PROPAGATE_2 10'b1000010111

//`define END_OF_PACKET_1 10'b1011101000
//`define END_OF_PACKET_2 10'b0100010111

//`define START_OF_PACKET_1 10'b1101101000
//`define START_OF_PACKET_2 10'b0010010111

//`define CARRIER_EXTEND_1 10'b1110101000
//`define CARRIER_EXTEND_2 10'b0001010111

//`define IDLE_1  10'b0011111010
//`define IDLE_2 10'b1100000101
//`define IDLE_3 10'b1010010110
//`define IDLE_4 10'b1010010110
//`define IDLE_5 10'b0110110101
//`define IDLE_6 10'b1001000101

//`define LP_IDLE_1  10'b0011111010
//`define LP_IDLE_2 10'b1100000101
//`define LP_IDLE_3 10'b0110011010
//`define LP_IDLE_4 10'b0110011010
//`define LP_IDLE_5 10'b0101101101
//`define LP_IDLE_6 10'b0101100010

//`define K28_5_N 10'b0011111010  
//`define K28_5_P 10'b1100000101

//`define D21_5 10'b1010101010

//`define D6_5 10'b0110011010 

//`define D5_6 10'b1010010110 

//`define D26_4_N 10'b0101101101 
//`define D26_4_P 10'b0101100010

//`define D16_2_N 10'b0110110101
//`define D16_2_P 10'b1001000101

`define K28_5 8'hBC
`define K27_7 8'hFB
`define K30_7 8'hFE
`define K23_7 8'hF7
`define K29_7 8'hFD
`define D21_5 8'hB5
`define D2_2 8'h42
`define D5_6 8'hC5
`define D16_2 8'h50
`define D0_0 8'h00

`define K28_5_10b_n 10'b0011111010
`define K28_5_10b_p 10'b1100000101

`define D21_5_10b_n 10'b1010101010
`define D21_5_10b_p 10'b1010101010

`define D2_2_10b_n 10'b1011010101
`define D2_2_10b_p 10'b0100100101

`define D5_6_10b_n 10'b1010010110
`define D5_6_10b_p 10'b1010010110

`define D16_2_10b_n 10'b0110110101
`define D16_2_10b_p 10'b1001000101

`define D6_5_10b_n 10'b0110011010
`define D6_5_10b_p 10'b0110011010

`define D26_4_10b_n 10'b0101101101
`define D26_4_10b_p 10'b0101100010

`define K27_7_10b_n 10'b1101101000
`define K27_7_10b_p 10'b0010010111




